`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: DD2 course 
// Engineer: Omar Shaalan
// ID: 900193887


//////////////////////////////////////////////////////////////////////////////////


module HA(sout,cout,a,b);
  output sout,cout;
  input a,b;
  assign sout=a^b;
  assign cout=(a&b);
endmodule
